reg rst_r;


wire clk100mhz;
wire locked, locked100;

wire rst_n;

wire rst0;


reg rst_x;

wire HDMI_CFG_READY;

assign rst0 = rst_r & locked & locked100;
assign rst = HDMI_CFG_READY & rst0;

assign clk = clk100mhz;


reg [17:0] resetcounter;

initial begin
   resetcounter <= 0;
   rst_r <= 0;
   rst_x <= 0;
end

// reset delay   
always @(posedge sys_clk_in)
  if (~rst_r) begin
     resetcounter <= resetcounter + 1;
     if (resetcounter[17]) rst_r <= 1;
  end

   always @(posedge sys_clk_in) begin
      rst_x <= rst_n;
   end



assign HDMI_I2S0  = 1'b z;
assign HDMI_MCLK  = 1'b z;
assign HDMI_LRCLK = 1'b z;
assign HDMI_SCLK  = 1'b z;
altera_pll# (
 .fractional_vco_multiplier("false"),
 .reference_clock_frequency("50 MHz"),
 .operation_mode("direct"),
 .number_of_clocks(1),
 .output_clock_frequency0("150 MHz"),
 .phase_shift0("0 ps"),
 .duty_cycle0(50),    
 .pll_type("General"),
 .pll_subtype("General")
)PLL2(
 .rst   (~rst_r),
 .outclk(clk100mhz),
 .locked(locked100),
 .refclk(sys_clk_in)
);

I2C_HDMI_Config #(
  .CLK_Freq (50000000),
  .I2C_Freq (20000) 
  )

  I2C_HDMI_Config (
  .iCLK        (sys_clk_in),
  .iRST_N      (rst0),
  .I2C_SCLK    (HDMI_I2C_SCL),
  .I2C_SDAT    (HDMI_I2C_SDA),
  .HDMI_TX_INT (HDMI_TX_INT),
  .READY       (HDMI_CFG_READY)
);

   wire [7:0] pseudoled;
   wire [7:0] pseudoled1;

   assign LED[0] = locked100;
   assign LED[1] = locked;
   assign LED[2] = HDMI_CFG_READY;
   
   
  
   ledwriter ledwr1 (.clk(clk),
                     .rst(rst),
                     
                     .LED({LED[7:3],pseudoled1[2:0]}),
                     
                     .addr_b(ram_addr_in_b),
                     .data_b_in(ram_data_out_b),
                     .data_b_we(ram_we_out));


`ifdef VGA4BIT

wire       clk25mhz;
   

// generate a PLL instance: 50MHz ref clock from the board,
// 25MHz output for VGA, 100MHz output for the rest of the SoC 
altera_pll# (
 .fractional_vco_multiplier("false"),
 .reference_clock_frequency("50 MHz"),
 .operation_mode("direct"),
 .number_of_clocks(1),
 .output_clock_frequency0("25 MHz"),
 .phase_shift0("0 ps"),
 .duty_cycle0(50),    
 .pll_type("General"),
 .pll_subtype("General")
)PLL1(
 .rst   (~rst_r),
 .outclk(clk25mhz),
 .locked(locked),
 .refclk(sys_clk_in)
);

   
wire vga_clsrq;

wire vga_clsack;

wire [19:0] vmem_in_addr;

wire [7:0] vmem_in_data;
wire [7:0] vmem_p1_out_data;

wire vmem_we;
wire vmem_re;

wire vmem_select;

wire vmem_bufswap;
wire vga_scan;


wire                    [3:0]   rgb;
assign HDMI_TX_CLK = clk25mhz;
   
assign HDMI_TX_D[23:16] = {rgb, 4'b0};
assign HDMI_TX_D[15:8] = {rgb, 4'b0};
assign HDMI_TX_D[7:0] = {rgb, 4'b0};

vgatopgfx vga1(.clk(clk),
               .rst(rst),

               .clk25mhz(clk25mhz),
               
	       .hsync(HDMI_TX_HS),
	       .vsync(HDMI_TX_VS),
	       .rgb(rgb),
               .dataenable(HDMI_TX_DE),
               
               .clsrq(vga_clsrq),
               .clsack(vga_clsack),
               .vmem_in_addr(vmem_in_addr),
               .vmem_in_data(vmem_in_data),
               .vmem_we(vmem_we),
               .vmem_re(vmem_re),
               .vmem_p1_out_data(vmem_p1_out_data),

               .bufswap(vmem_bufswap),
               .vga_scan(vga_scan)
               );

`endif //  `ifdef VGA4BIT

`ifdef BIGMEM
   
wire clk_vga; // 148.5MHz generated by the soc_system PLL
   
wire  [27:0] vbuf_address;
wire   [7:0] vbuf_burstcount;
wire         vbuf_waitrequest;
wire [127:0] vbuf_readdata;
wire         vbuf_readdatavalid;
wire         vbuf_read;
wire [127:0] vbuf_writedata;
wire  [15:0] vbuf_byteenable;
wire         vbuf_write;
   assign vbuf_write = 0;
   assign vbuf_writedata = 0;
   assign vbuf_byteenable = 0;
   

   
   wire [28:0] ram1_address;
   wire [7:0] ram1_burstcount;
   wire    ram1_waitrequest;

   wire [63:0] ram1_readdata;
   wire     ram1_readdatavalid;
   wire     ram1_read;
   wire [63:0] ram1_writedata;
   wire [7:0] ram1_byteenable;
   wire     ram1_write;


   wire [1:0] vga_bufid;
   wire       vga_scan;
   
   wire [23:0] rgb;
   assign HDMI_TX_CLK = clk_vga;
   
   assign HDMI_TX_D = rgb;

vga1080p vga    (.clk(clk),
		 .clk_vga(clk_vga),
		 .rst(rst),
		 .bufid(vga_bufid),
		 .vbuf_address(vbuf_address),
		 .vbuf_burstcount(vbuf_burstcount),
		 .vbuf_readdata(vbuf_readdata),
		 .vbuf_readdatavalid(vbuf_readdatavalid),
		 .vbuf_read(vbuf_read),
		 .scan(vga_scan),
		 
		 .LED(pseudoled),
		 
		 .hsync(HDMI_TX_HS),
		 .vsync(HDMI_TX_VS),
		 .rgb(rgb),
		 .dataenable(HDMI_TX_DE));

soc_system u0  (
		.clk_clk                             (sys_clk_in),                             //                    clk.clk
		.ddr3_clk_clk                        (clk_vga),

		.pll_locked_export                          (locked),

		.ddr3_hps_f2h_sdram0_clock_clk          (clk),          // hps_0_f2h_sdram0_clock.clk

		.ddr3_hps_f2h_sdram1_data_address       (ram1_address),       //  hps_0_f2h_sdram0_data.address
		.ddr3_hps_f2h_sdram1_data_burstcount    (ram1_burstcount),    //                       .burstcount
		.ddr3_hps_f2h_sdram1_data_waitrequest   (ram1_waitrequest),   //                       .waitrequest
		.ddr3_hps_f2h_sdram1_data_readdata      (ram1_readdata),      //                       .readdata
		.ddr3_hps_f2h_sdram1_data_readdatavalid (ram1_readdatavalid), //                       .readdatavalid
		.ddr3_hps_f2h_sdram1_data_read          (ram1_read),          //                       .read
		.ddr3_hps_f2h_sdram1_data_writedata     (ram1_writedata),     //                       .writedata
		.ddr3_hps_f2h_sdram1_data_byteenable    (ram1_byteenable),    //                       .byteenable
		.ddr3_hps_f2h_sdram1_data_write         (ram1_write),         //                       .write

		.ddr3_hps_f2h_sdram0_data_address       (vbuf_address),       //  hps_0_f2h_sdram1_data.address
		.ddr3_hps_f2h_sdram0_data_burstcount    (vbuf_burstcount),    //                       .burstcount
		.ddr3_hps_f2h_sdram0_data_waitrequest   (vbuf_waitrequest),   //                       .waitrequest
		.ddr3_hps_f2h_sdram0_data_readdata      (vbuf_readdata),      //                       .readdata
		.ddr3_hps_f2h_sdram0_data_readdatavalid (vbuf_readdatavalid), //                       .readdatavalid
		.ddr3_hps_f2h_sdram0_data_read          (vbuf_read),          //                       .read
		.ddr3_hps_f2h_sdram0_data_writedata     (vbuf_writedata),     //                       .writedata
		.ddr3_hps_f2h_sdram0_data_byteenable    (vbuf_byteenable),    //                       .byteenable
		.ddr3_hps_f2h_sdram0_data_write         (vbuf_write),         //                       .write

		// A second 65-bit port
		.ddr3_hps_f2h_sdram2_data_address       (0),       //  hps_0_f2h_sdram1_data.address
		.ddr3_hps_f2h_sdram2_data_burstcount    (0),    //                       .burstcount
		.ddr3_hps_f2h_sdram2_data_waitrequest   (),   //                       .waitrequest
		.ddr3_hps_f2h_sdram2_data_readdata      (),      //                       .readdata
		.ddr3_hps_f2h_sdram2_data_readdatavalid (), //                       .readdatavalid
		.ddr3_hps_f2h_sdram2_data_read          (0),          //                       .read
		.ddr3_hps_f2h_sdram2_data_writedata     (0),     //                       .writedata
		.ddr3_hps_f2h_sdram2_data_byteenable    (0),    //                       .byteenable
		.ddr3_hps_f2h_sdram2_data_write         (0),         //                       .write

		//HPS ddr3
		.memory_mem_a                          ( HPS_DDR3_ADDR),                       //                memory.mem_a
		.memory_mem_ba                         ( HPS_DDR3_BA),                         //                .mem_ba
		.memory_mem_ck                         ( HPS_DDR3_CK_P),                       //                .mem_ck
		.memory_mem_ck_n                       ( HPS_DDR3_CK_N),                       //                .mem_ck_n
		.memory_mem_cke                        ( HPS_DDR3_CKE),                        //                .mem_cke
		.memory_mem_cs_n                       ( HPS_DDR3_CS_N),                       //                .mem_cs_n
		.memory_mem_ras_n                      ( HPS_DDR3_RAS_N),                      //                .mem_ras_n
		.memory_mem_cas_n                      ( HPS_DDR3_CAS_N),                      //                .mem_cas_n
		.memory_mem_we_n                       ( HPS_DDR3_WE_N),                       //                .mem_we_n
		.memory_mem_reset_n                    ( HPS_DDR3_RESET_N),                    //                .mem_reset_n
		.memory_mem_dq                         ( HPS_DDR3_DQ),                         //                .mem_dq
		.memory_mem_dqs                        ( HPS_DDR3_DQS_P),                      //                .mem_dqs
		.memory_mem_dqs_n                      ( HPS_DDR3_DQS_N),                      //                .mem_dqs_n
		.memory_mem_odt                        ( HPS_DDR3_ODT),                        //                .mem_odt
		.memory_mem_dm                         ( HPS_DDR3_DM),                         //                .mem_dm
		.memory_oct_rzqin                      ( HPS_DDR3_RZQ),                        //                .oct_rzqin
		//HPS SPI
		.hps_io_hps_io_spim1_inst_CLK(HPS_SPIM_CLK),           //                               .hps_io_spim1_inst_CLK
		.hps_io_hps_io_spim1_inst_MOSI(HPS_SPIM_MOSI),         //                               .hps_io_spim1_inst_MOSI
		.hps_io_hps_io_spim1_inst_MISO(HPS_SPIM_MISO),         //                               .hps_io_spim1_inst_MISO
		.hps_io_hps_io_spim1_inst_SS0(HPS_SPIM_SS),            //                               .hps_io_spim1_inst_SS0

                //HPS SD card
               .hps_io_hps_io_sdio_inst_CMD(HPS_SD_CMD),              //                               .hps_io_sdio_inst_CMD
               .hps_io_hps_io_sdio_inst_D0(HPS_SD_DATA[0]),           //                               .hps_io_sdio_inst_D0
               .hps_io_hps_io_sdio_inst_D1(HPS_SD_DATA[1]),           //                               .hps_io_sdio_inst_D1
               .hps_io_hps_io_sdio_inst_CLK(HPS_SD_CLK),              //                               .hps_io_sdio_inst_CLK
               .hps_io_hps_io_sdio_inst_D2(HPS_SD_DATA[2]),           //                               .hps_io_sdio_inst_D2
               .hps_io_hps_io_sdio_inst_D3(HPS_SD_DATA[3]),           //                               .hps_io_sdio_inst_D3
               //HPS UART
               .hps_io_hps_io_uart0_inst_RX(HPS_UART_RX),             //                               .hps_io_uart0_inst_RX
               .hps_io_hps_io_uart0_inst_TX(HPS_UART_TX),             //                               .hps_io_uart0_inst_TX
               //HPS I2C1
               .hps_io_hps_io_i2c0_inst_SDA(HPS_I2C0_SDAT),           //                               .hps_io_i2c0_inst_SDA
               .hps_io_hps_io_i2c0_inst_SCL(HPS_I2C0_SCLK),           //                               .hps_io_i2c0_inst_SCL
               //HPS I2C2
               .hps_io_hps_io_i2c1_inst_SDA(HPS_I2C1_SDAT),           //                               .hps_io_i2c1_inst_SDA
               .hps_io_hps_io_i2c1_inst_SCL(HPS_I2C1_SCLK)            //                               .hps_io_i2c1_inst_SCL

		);
   

`endif
